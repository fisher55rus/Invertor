* C:\Workspace_git\Magistr\Shevtsov\Invertor\Orcad\3_Limit\Limit.sch

* Schematics Version 9.2
* Mon Feb 18 18:54:14 2019



** Analysis setup **
.tran 0ns 60m 0 1.57u SKIPBP
.LIB "C:\Workspace_git\Magistr\Shevtsov\Invertor\Orcad\2_Sinus_generator\Sinus_generator.lib"


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "Limit.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
