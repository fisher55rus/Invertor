* D:\GIT\MAI\Invertor\Orcad\2_Sinus_generator\SG_prec.sch

* Schematics Version 9.2
* Fri Apr 12 18:38:15 2019



** Analysis setup **
.tran 0ns 100m 0 1.57u SKIPBP
.LIB "D:\GIT\MAI\Invertor\Orcad\2_Sinus_generator\Sinus_generator.lib"


* From [PSPICE NETLIST] section of d:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "D:\Program Files\Orcad\PSpice\UserLib\OPA_2.lib"
.lib "D:\Program Files\Orcad\PSpice\UserLib\MyLib.lib"
.lib "nom.lib"

.INC "SG_prec.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
