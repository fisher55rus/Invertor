* C:\Program Files\Orcad\work\Magistr2\1STK.sch

* Schematics Version 9.2
* Mon Feb 11 19:26:49 2019



** Analysis setup **
.tran 0ns 200us 0 1.57u SKIPBP
.OPTIONS ABSTOL=1uA
.OPTIONS ITL4=60
.LIB "C:\Program Files\Orcad\work\Magistr2\1STK.lib"


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "1STK.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
