* D:\GIT\MAI\Invertor\Orcad\11_constant_current_transform\trash\Schematic2.sch

* Schematics Version 9.2
* Sun Apr 21 20:31:24 2019


.PARAM         Ep=27 Rvar=5 

** Analysis setup **
.tran 0ns 50ms 0 1.57u SKIPBP
.OPTIONS ABSTOL=1uA
.OPTIONS ITL4=60
.OPTIONS RELTOL=0.01
.LIB "D:\GIT\MAI\Invertor\Orcad\Test_Var\Schematic2.lib"


* From [PSPICE NETLIST] section of d:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "D:\Program Files\Orcad\PSpice\UserLib\OPA_2.lib"
.lib "D:\Program Files\Orcad\PSpice\UserLib\MyLib.lib"
.lib "nom.lib"

.INC "Schematic2.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
