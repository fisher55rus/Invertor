* D:\GIT\MAI\Invertor\Orcad\1_Power_cascade\1STK.sch

* Schematics Version 9.2
* Wed Apr 10 21:45:11 2019



** Analysis setup **
.tran 0ns 200u 0 1.57u SKIPBP
.OPTIONS ABSTOL=1uA
.OPTIONS ITL4=60
.LIB "D:\GIT\MAI\Invertor\Orcad\1_Power_cascade\1STK.lib"


* From [PSPICE NETLIST] section of d:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "D:\Program Files\Orcad\PSpice\UserLib\OPA_2.lib"
.lib "D:\Program Files\Orcad\PSpice\UserLib\MyLib.lib"
.lib "nom.lib"

.INC "1STK.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
