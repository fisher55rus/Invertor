* D:\GIT\MAI\Invertor\Orcad\10_DC_sweep_27v_10-500ohm\test.sch

* Schematics Version 9.2
* Sun Apr 21 19:40:55 2019


.PARAM         Rn=5 

** Analysis setup **
.tran 0ns 5ms 2.5ms 1.57u SKIPBP
.four 400 99 V([V_sence])
.STEP  PARAM Rn LIST 
+ 5, 50, 100, 150, 200, 250, 300, 350, 400, 450, 500
.LIB "D:\GIT\MAI\Invertor\Orcad\1_Power_cascade\1STK.lib"


* From [PSPICE NETLIST] section of d:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "D:\Program Files\Orcad\PSpice\UserLib\OPA_2.lib"
.lib "D:\Program Files\Orcad\PSpice\UserLib\MyLib.lib"
.lib "nom.lib"

.INC "test.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
