* C:\Workspace_git\Magistr\Shevtsov\Invertor\Orcad\7_full3\1STK.sch

* Schematics Version 9.2
* Mon Feb 25 19:02:37 2019



** Analysis setup **
.tran 0ns 10m 0 1.57u SKIPBP
.OPTIONS ABSTOL=1uA
.OPTIONS ITL4=60
.LIB "C:\Workspace_git\Magistr\Shevtsov\Invertor\Orcad\6_full2\1STK.lib"


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "C:\Program Files\Orcad\PSpice\UserLib\Mylib.lib"
.lib "nom.lib"
.inc "C:\Program Files\Orcad\PSpice\UserLib\Mylib.lib"

.INC "1STK.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
