* D:\GIT\MAI\Invertor\Orcad\16_Driver_with_pervi4ka\Schematic2.sch

* Schematics Version 9.2
* Mon Mar 11 18:55:31 2019



** Analysis setup **
.tran 0ns 200u 0 0.1u SKIPBP
.LIB "D:\GIT\MAI\Invertor\Orcad\15_Driver_with_stab\Schematic2.lib"


* From [PSPICE NETLIST] section of d:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "D:\Program Files\Orcad\PSpice\UserLib\OPA_2.lib"
.lib "D:\Program Files\Orcad\PSpice\UserLib\MyLib.lib"
.lib "nom.lib"

.INC "Schematic2.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
