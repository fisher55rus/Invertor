* D:\GIT\MAI\Invertor\Orcad\14_Driver\Schematic2.sch

* Schematics Version 9.2
* Mon Mar 11 17:57:56 2019



** Analysis setup **
.tran 0ns 200u 0 0.1u SKIPBP


* From [PSPICE NETLIST] section of d:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "D:\Program Files\Orcad\PSpice\UserLib\OPA_2.lib"
.lib "D:\Program Files\Orcad\PSpice\UserLib\MyLib.lib"
.lib "nom.lib"

.INC "Schematic2.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
