* D:\GIT\MAI\Invertor\Orcad\6_full2\test.sch

* Schematics Version 9.2
* Sat Apr 13 11:15:39 2019



** Analysis setup **
.tran 0ns 10m 0 1.57u SKIPBP
.LIB "D:\GIT\MAI\Invertor\Orcad\1_Power_cascade\1STK.lib"


* From [PSPICE NETLIST] section of d:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "D:\Program Files\Orcad\PSpice\UserLib\OPA_2.lib"
.lib "D:\Program Files\Orcad\PSpice\UserLib\MyLib.lib"
.lib "nom.lib"

.INC "test.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
